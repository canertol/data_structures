module instmem (a,rd,rd1512);
input [31:0] a;
output [31:0] rd;
output [15:12] rd1512;

reg [31:0] inst[63:0];

initial begin
 inst[4]=32'b11100010100000000010000000000111;  // r2=5 ADD R2, R0, #5
 inst[8]=32'b11100010100000000011000000001100;  // r3=12 ADD R3, R0, #12
 inst[12]=32'b11100010010000110111000000001001; // r7=3 SUB R7, R3, #9
 inst[16]=32'b11100001100001110100000000000010; // r4= 3or5 = 7 ORR R4, R7, R2
 inst[20]=32'b11100000000000110101000000000100; // r5=12and7 = 4 AND R5, R3, R4
 inst[24]=32'b11100000100001010101000000000100; // r5=4+7=11  ADD R5, R5, R4
 inst[28]=32'b11100101100000110111000001010100; // mem[12+84]=3 STR R7, [R3, #84]
 inst[32]=32'b11100101100100000010000001100000; // r2=mem[96]=3 LDR R2, [R0, #96]
 inst[36]=32'b11100001010101000000000000000010; // cmp r4 r2
 inst[40]=32'b11100001101000000010000010100011; //lsr r2 r3 1
 inst[44]=32'b11100001101000000010000010000011; //lsl r2 r3 1
 end
assign rd= inst[a[31:0]];
assign rd1512=inst[a[31:0]][15:12];

endmodule