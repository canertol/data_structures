module INST_MEM (A,RD);
input [31:0] A;
output [31:0] RD;

reg [31:0] INST[92:0];

initial begin
 INST[0]  = 32'b1110_000_0010_0_1111_0000_0000_0000_1111; //	    SUB R0, R15, R15 	; R0 = 0
 INST[4]  = 32'b1110_001_0100_0_0000_0010_0000_0000_0101; // 		 ADD R2, R0, #5 		; R2 = 5
 INST[8]  = 32'b1110_001_0100_0_0000_0011_0000_0000_1100; // 		 ADD R3, R0, #12		; R3 = 12
 INST[12] = 32'b1110_001_0010_0_0011_0111_0000_0000_1001; // 		 SUB R7, R3, #9 		; R7 = 3
 INST[16] = 32'b1110_000_1100_0_0111_0100_0000_0000_0010; // 		 ORR R4, R7, R2 		; R4 = 3 OR 5 = 7
 INST[20] = 32'b1110_000_0000_0_0011_0101_0000_0000_0100; // 		 AND R5, R3, R4 		; R5 = 12 AND 7 = 4
 INST[24] = 32'b1110_000_0100_0_0101_0101_0000_0000_0100; // 		 ADD R5, R5, R4 		; R5 = 4 + 7 = 11
 INST[28] = 32'b1110_000_0010_1_0101_1000_0000_0000_0111; // 		 SUB R8, R5, R7 		; R8 = 11 - 3 = 8
 
 INST[32] = 32'b1110_010_1100_0_0000_0010_1000_0000_0000; //		 STR  R2, R8 	      ; R2 = R8 = 7
 INST[36] = 32'b1110_010_1100_1_0000_0010_1000_0000_0000; //		 LDR  R2, R8 	      ; R2 = R8 = 7
/*
 INST[36] = 32'b1110_000_0010_1_0011_1000_0000_0000_0100; // 		 SUBS R8, R3, R4 		; R8 = 12 - 7 = 5
 INST[40] = 32'b1110_000_1101_0_0000_0010_0000_1010_0011; //		 LSR  R2, R3, #1
 INST[44] = 32'b1110_001_0100_0_0000_0101_0000_0000_0000; // 		 ADD R5, R0, #0 		; should be skipped
 INST[48] = 32'b1110_000_0010_1_0111_1000_0000_0000_0010; //       SUBS R8, R7, R2 		; R8 = 3 - 5 = -2, set Flags
 INST[52] = 32'b1011_001_0100_0_0101_0111_0000_0000_0001; //		 ADDLT R7, R5, #1 	; R7 = 11 + 1 = 12
 INST[56] = 32'b1110_000_0010_0_0111_0111_0000_0000_0010; // 		 SUB R7, R7, R2 		; R7 = 12 - 5 = 7
 INST[60] = 32'b1110_010_1100_0_0011_0111_0000_0101_0100; //		 STR R7, [R3, #84] 	; mem[12+84] = 7
 INST[64] = 32'b1110_010_1100_1_0000_0010_0000_0110_0000; //		 LDR R2, [R0, #96] 	; R2 = mem[96] = 7
 INST[68] = 32'b1110_000_0100_0_1111_1111_0000_0000_0000; //		 ADD R15, R15, R0 	; PC = PC+8 (skips next)
 INST[72] = 32'b1110_001_0100_0_0000_0010_0000_0000_0001; //		 ADD R2, R0, #14 		; shouldn't happen
 INST[76] = 32'b1110_000_1010_1_0100_0000_0000_0000_0010; 			 // 	    CMP R4, R2
 INST[80] = 32'b1110_001_0100_0_0000_0010_0000_0000_0001; //		 ADD R2, R0, #13 		; shouldn't happen
 INST[84] = 32'b1110_001_0100_0_0000_0010_0000_0000_0001; //		 ADD R2, R0, #10 		; shouldn't happen
 INST[88] = 32'b1110_010_1100_0_0000_0010_0000_0101_0100;  //       STR R2, [R0, #100]  ; mem[100] = 7
 INST[92] = 32'b1110_000_1101_0_000_0001_0000_0100_00011; 			 //		 lsl r2 r3 1
 */
end 

assign RD = INST[A];

endmodule