module register_file  #(parameter, W = 3)(
       clk, 
       WD3, WE3, rst
       A1, A2, A3, 
       RD1, RD2);
  
       // inputs
       input clk;
       input [W:0] data_in;
       input [1:0] A1, A2, A3;
       input WE3, rst;
       // outputs
       output reg [W:0] RD1, RD2;
  
  
  
  
  
  
endmodule
