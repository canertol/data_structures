module register_file  #(parameter, W = 3)(data_in, data_out1, data_out2)

endmodule
