module IDM(A, WD, clk, WE, out); 
 input [7:0] WD;                    
 input[7:0] A;
 input clk, WE;
 output [15:0] out;
 reg [15:0] data[63:0]; // 2^6 memory slots
 
 initial begin
 // INSTRUCTION PART /////////////////////////////////////
	 data[0]<=16'b10_001_110_00001010; // BLD #10
	 data[1]<=16'b10_000_110_00011101; // BUN #29
	 data[2]<=16'b10_001_110_00101000; // BLD #40
	 data[3]<=16'b11_000_01000000000; //finish

 // Subroutine 1 - Memory Instructions	 
	 data[10]<=16'b11_000_010_00000001; // LDD R2, #1			; R2 = 1
	 data[11]<=16'b11_000_011_00000100; // LDD R3, #4			; R3 = 4
	 data[12]<=16'b11_010_011_00110111;	// STD R3, [#55]		; M[55] = 4
	 data[13]<=16'b11_001_010_00110111;	// LDM R2,[#55]		; R2 = 4
	 data[14]<=16'b11_000_010_00000110; // LDD R2, #6			; R2 = 6
	 data[15]<=16'b10_001_110_00000001; // BLD #1
	 
	  // DATA PART /////////////////////////////////////
	 data[16]<=4'h00_01;
	 data[17]<=4'h00_02;
	 data[18]<=4'h00_03;
	 data[19]<=4'h00_04;
	 data[20]<=4'h00_05;
	 data[21]<=4'h00_06;
	 data[22]<=4'h00_07;
	 data[23]<=4'h00_08;
	 data[24]<=4'h00_09;
	 data[25]<=4'h00_0A;
	 data[26]<=4'h00_0B;
	 data[27]<=4'h00_0C;
	 data[28]<=4'h00_0D;	 
	 /////////////////////////////////////
	 
 // Subroutine 2 - Arithmetic & Logic Instructions	 
	 data[29]<=16'b00_000_001_010_011_00; // ADD R1, R2, R3   ; R1 = 6 + 4 = 10
	 data[30]<=16'b00_001_100_001_011_00; // SUB R4, R1, R3	 ; R4 = 10 - 4 = 6
	 data[31]<=16'b00_010_010_011_10000;  // ADDI R2,R3,[#16]  ; R2 = 6 + 1 = 7 =10 *************
	 data[32]<=16'b00_011_000_010_10000;  // SUBI R0,R2,[#16]  ; R0 = 7- 1 = 6=4************
	 data[33]<=16'b00_100_000_000_010_00; // AND	R0,R0,R2		 ; R0 = 6 & 7 = 6 =0
	 data[34]<=16'b00_101_010_011_010_00; // ORR R2,R3,R2  	 ; R2 = 6 | 7 = 7 = 14
	 data[35]<=16'b00_110_000_010_001_00; // XOR R0,R2,R1		 ; R0 = 7 ^ 10 = 13 = 4
	 data[36]<=16'b00_111_000_000_000_00; // CLR R0				 ; R0 = 0
	 data[37]<=16'b10_100_110_00011101;   // BNE #2
	 data[38]<=16'b10_011_110_00000010;   // BEQ #2

 // Subroutine 3 - Shift Instructions
	 data[40]<=16'b01_000_001_001_00000;  // ROL R1				 ; R1 = 20
	 data[41]<=16'b01_001_010_010_00000;  // ROR R2				 ;	R2 = 8'b00000111
	 data[42]<=16'b01_001_010_010_00000;  // ROR R2				 ;	R2 = 8'b10000011
	 data[43]<=16'b01_010_100_100_00000;  // LSL R4				 ; R4 = 12
	 data[44]<=16'b01_011_010_010_00000;  // ASR R2				 ; R2 = 8'b11000001
	 data[45]<=16'b01_100_010_010_00000;  // LSR R2				 ; R2 = 8'b01100000
	 data[46]<=16'b10_001_110_00000011;   // BLD #3
	


	
 end
 
 always @(posedge clk)begin
  if(WE) data[A[7:0]]<= WD;
 end
 
 assign out = data[A[7:0]];
endmodule
 