module controller(
                CLK, RST,
                AccRight, AccParallel, // Acc register control
                OP, ASrc, BSrc,  // ALU Controllers
                Stat, NFlag,    // Status bits
                INST // Instruction
              );





endmodule
